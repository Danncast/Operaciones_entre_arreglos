
library ieee;
use ieee.std_logic_1164.all;

--Entity
Entity Comparator is
	generic ( n: integer :=7);--<-- nbits
	Port(
		Addr , B: in std_logic_vector(n-1 downto 0);
		AmenorB, AmayorB, AigualB: out std_logic);
end Comparator;

--Architecture
Architecture solve of Comparator is
	-- Signals,Constants,Variables,Components
	Begin
		AmenorB<='1' when Addr<B else '0';
		AmayorB<='1' when Addr>B else '0';
		AigualB<='1' when Addr=B else '0';
end solve;